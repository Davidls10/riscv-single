module instruction_memory(input wire [31:0] pc,
                          output reg [31:0] instr);

    /*
    L7: lw x6, -4(x9)        I   111111111100 01001 010 00110 0000011
        sw x6, 8(x9)         S   0000000 00110 01001 010 01000 0100011
        or x4, x5, x6        R   0000000 00110 00101 110 00100 0110011
        addi x4, x4, 2       I   000000000010 00100 000 00100 0010011
        and x4, x4, x6       R   0000000 00110 00100 111 00100 0110011
        beq x4, x4, L7       B   1111111 00100 00100 000 01101 1100011
    */

    always @* begin
        case(pc)
            32'h0000: instr = 32'b11111111110001001010001100000011;
            32'h0004: instr = 32'b00000000011001001010010000100011;
            32'h0008: instr = 32'b00000000011000101110001000110011;
            32'h000c: instr = 32'b00000000001000100000001000010011;
            32'h0010: instr = 32'b00000000011000100111001000110011;
            32'h0014: instr = 32'b11111110010000100000011011100011;
        endcase
    end
    
endmodule