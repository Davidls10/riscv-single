module instruction_memory(input wire [15:0] pc,
                          output wire [31:0] instr);

    /*
    L7: lw x6, -4(x9)        I   111111111100 01001 010 00110 0000011
        sw x6, 8(x9)         S   0000000 00110 01001 010 01000 0100011
        or x4, x5, x6        R   0000000 00110 00101 110 00100 0110011 
        beq x4, x4, L7       B   1111111 00100 00100 000 10101 1100011
    */

    always @* begin
        case(pc)
            16'h00: instr = 32'b11111111110001001010001100000011;
            16'h04: instr = 32'b00000000011001001010010000100011;
            16'h08: instr = 32'b00000000011000101110001000110011;
            16'h0c: instr = 32'b11111110010000100000101011100011;
        endcase
    end
    
endmodule