module decoder#(parameter N = 8)
               (output wire )

    
endmodule